package ov5640_1080p30_pkg;

parameter bit [36 : 0][23 : 0] MODE_ROM = {
  24'h3008_02,
  24'h501f_03,
  24'h4300_00,
  24'h370c_03,
  24'h3709_52,
  24'h3708_64,
  24'h3612_59,
  24'h3618_00,
  24'h4837_14,
  24'h3821_00,
  24'h3815_11,
  24'h3814_11,
  24'h380f_60,
  24'h380e_04,
  24'h380d_c4,
  24'h380c_09,
  24'h380b_38,
  24'h380a_04,
  24'h3809_80,
  24'h3808_07,
  24'h3813_0c,
  24'h3812_00,
  24'h3811_10,
  24'h3810_00,
  24'h3807_f9,
  24'h3806_05,
  24'h3805_ef,
  24'h3804_08,
  24'h3803_aa,
  24'h3802_01,
  24'h3801_50,
  24'h3800_01,
  24'h3034_1a,
  24'h3108_01,
  24'h3037_15,
  24'h3036_54,
  24'h3035_11 };
  
parameter int TOTAL_MODE_OPS = 37;

endpackage
