package ov5640_init_pkg;

parameter bit [63 : 0][23 : 0] INIT_ROM = {
  24'h5001_00,
  24'h5000_00,
  24'h3824_01,
  24'h460c_20,
  24'h460b_35,
  24'h440e_00,
  24'h4407_04,
  24'h4818_01,
  24'h4713_03,
  24'h501f_01,
  24'h4300_6f,
  24'h302e_08,
  24'h4800_14,
  24'h300e_45,
  24'h3820_46,
  24'h503d_00,
  24'h3c0b_40,
  24'h3c0a_9c,
  24'h3c09_1c,
  24'h3c08_00,
  24'h3c07_08,
  24'h3c06_00,
  24'h3c05_98,
  24'h3c04_28,
  24'h3c01_34,
  24'h3622_01,
  24'h3634_44,
  24'h3636_06,
  24'h3635_13,
  24'h3a19_f8,
  24'h3a18_00,
  24'h3a13_43,
  24'h471c_50,
  24'h371b_20,
  24'h3620_52,
  24'h302d_60,
  24'h3601_33,
  24'h3600_37,
  24'h3731_02,
  24'h3901_0a,
  24'h3906_10,
  24'h3905_02,
  24'h3705_1a,
  24'h370b_60,
  24'h3717_01,
  24'h3715_78,
  24'h3703_5a,
  24'h3704_a0,
  24'h3621_e0,
  24'h3633_23,
  24'h3632_e2,
  24'h3631_0e,
  24'h3630_2e,
  24'h303b_19,
  24'h303d_10,
  24'h3108_01,
  24'h3037_11,
  24'h3036_38,
  24'h3035_11,
  24'h3034_18,
  24'h3018_00,
  24'h3017_00,
  24'h3103_03,
  24'h3008_42
};

parameter int TOTAL_INIT_OPS = 64;

endpackage
