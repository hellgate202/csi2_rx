package imx477_1080p30_pkg;

parameter bit [104 : 0][23 : 0] MODE_ROM = {
  24'h0100_01,
  24'h0341_6e,
  24'h0340_04,
  24'h0205_00,
  24'h0204_00,
  24'h0203_40,
  24'h0202_04,
  24'h0101_00,
  24'h3f57_6c,
  24'h3f56_01,
  24'h3f50_00,
  24'h3e37_00,
  24'h3e20_01,
  24'he04f_1f,
  24'he04e_00,
  24'he04d_7f,
  24'he04c_00,
  24'h0819_3f,
  24'h0818_00,
  24'h0817_27,
  24'h0816_01,
  24'h0815_4f,
  24'h0814_00,
  24'h0813_57,
  24'h0812_00,
  24'h0811_5f,
  24'h0810_00,
  24'h080f_77,
  24'h080e_00,
  24'h080d_4f,
  24'h080c_00,
  24'h080b_7f,
  24'h080a_00,
  24'h0823_00,
  24'h0822_00,
  24'h0821_08,
  24'h0820_07,
  24'h0310_01,
  24'h030f_7d,
  24'h030e_00,
  24'h030d_02,
  24'h030b_02,
  24'h0309_0a,
  24'h0307_5e,
  24'h0306_01,
  24'h0305_04,
  24'h0303_02,
  24'h0301_05,
  24'h034f_38,
  24'h034e_04,
  24'h034d_ec,
  24'h034c_07,
  24'h040f_38,
  24'h040e_04,
  24'h040d_d8,
  24'h040c_0f,
  24'h040b_00,
  24'h040a_00,
  24'h0409_00,
  24'h0408_00,
  24'h0405_20,
  24'h0404_00,
  24'h0401_01,
  24'ha2b7_00,
  24'ha2a9_60,
  24'h9e9f_00,
  24'h9e9e_00,
  24'h9e9d_00,
  24'h9e9c_2f,
  24'h9e9b_2f,
  24'h9e9a_2f,
  24'h9305_00,
  24'h9304_00,
  24'h936d_5f,
  24'h936b_64,
  24'h9369_73,
  24'h7b53_01,
  24'h574b_00,
  24'h574a_00,
  24'h5749_ff,
  24'h5748_07,
  24'h3f0d_01,
  24'h3c02_a2,
  24'h3c01_03,
  24'h3c00_00,
  24'h3140_02,
  24'h0902_02,
  24'h0901_12,
  24'h0900_01,
  24'h0387_01,
  24'h0385_01,
  24'h0383_01,
  24'h0381_01,
  24'h0221_11,
  24'h0220_00,
  24'h034b_27,
  24'h034a_0a,
  24'h0349_d7,
  24'h0348_0f,
  24'h0347_b8,
  24'h0346_01,
  24'h0345_00,
  24'h0344_00,
  24'h0343_c4,
  24'h0342_5f
};
  
parameter int TOTAL_MODE_OPS = 105;

endpackage
