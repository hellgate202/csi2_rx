package csi2_err_bit_pos_pkg;

parameter bit [63 : 0][7 : 0] ROM_INIT = {
  5'h1F,
  5'h1F,
  5'h1F,
  5'h1F,
  5'h1F,
  5'h1F,
  5'h1F,
  5'h00,
  5'h1F,
  5'h1F,
  5'h1F,
  5'h01,
  5'h1F,
  5'h02,
  5'h03,
  5'h1F,
  5'h1F,
  5'h1F,
  5'h1F,
  5'h04,
  5'h1F,
  5'h05,
  5'h06,
  5'h1F,
  5'h1F,
  5'h07,
  5'h08,
  5'h1F,
  5'h09,
  5'h1F,
  5'h1F,
  5'h14,
  5'h1F,
  5'h1F,
  5'h1F,
  5'h0A,
  5'h1F,
  5'h0B,
  5'h0C,
  5'h1F,
  5'h1F,
  5'h0D,
  5'h0E,
  5'h1F,
  5'h0F,
  5'h1F,
  5'h1F,
  5'h15,
  5'h1F,
  5'h10,
  5'h11,
  5'h1F,
  5'h12,
  5'h1F,
  5'h1F,
  5'h16,
  5'h13,
  5'h1F,
  5'h1F,
  5'h17,
  5'h1F,
  5'h1F,
  5'h1F,
  5'h1F };

endpackage
