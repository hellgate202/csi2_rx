package imx477_init_pkg;

parameter bit [307 : 0][23 : 0] INIT_ROM = {
  24'hbcf1_02,
  24'h0350_00,
  24'h0114_01,
  24'h0113_0c,
  24'h0112_0c,
  24'hb35e_08,
  24'hb35c_00,
  24'hb21f_04,
  24'ha2b9_00,
  24'ha2ad_ff,
  24'ha257_00,
  24'ha24b_ff,
  24'ha1b9_00,
  24'ha1b5_50,
  24'ha1b3_0c,
  24'ha1ad_ff,
  24'ha157_00,
  24'ha155_02,
  24'ha153_50,
  24'ha151_0c,
  24'ha148_ff,
  24'h9fcd_0a,
  24'h9fcb_0a,
  24'h9fc9_0a,
  24'h9fae_09,
  24'h9fad_09,
  24'h9fac_09,
  24'h9fab_00,
  24'h9faa_00,
  24'h9fa9_00,
  24'h9fa8_1e,
  24'h9fa7_1e,
  24'h9fa6_1e,
  24'h9fa5_00,
  24'h9fa4_00,
  24'h9fa3_00,
  24'h9fa2_0f,
  24'h9fa1_0f,
  24'h9fa0_0f,
  24'h9f9f_00,
  24'h9f9e_00,
  24'h9f9d_00,
  24'h9f9c_2f,
  24'h9f9b_2f,
  24'h9f9a_2f,
  24'h9f99_00,
  24'h9f98_00,
  24'h9f97_00,
  24'h9f96_0f,
  24'h9f95_0f,
  24'h9f94_0f,
  24'h9f75_04,
  24'h9f73_32,
  24'h9f71_c8,
  24'h9f6b_00,
  24'h9f4d_5a,
  24'h9f47_42,
  24'h9f41_6b,
  24'h9f3b_2f,
  24'h9f29_50,
  24'h9f1d_31,
  24'h9f17_35,
  24'h9ecd_0a,
  24'h9ecb_0a,
  24'h9ec9_0a,
  24'h9eae_09,
  24'h9ead_09,
  24'h9eac_09,
  24'h9eab_00,
  24'h9eaa_00,
  24'h9ea9_00,
  24'h9ea8_3f,
  24'h9ea7_3f,
  24'h9ea6_3f,
  24'h9ea5_00,
  24'h9ea4_00,
  24'h9ea3_00,
  24'h9ea2_0f,
  24'h9ea1_0f,
  24'h9ea0_0f,
  24'h9e99_00,
  24'h9e98_00,
  24'h9e97_00,
  24'h9e96_0f,
  24'h9e95_0f,
  24'h9e94_0f,
  24'h9e75_04,
  24'h9e73_32,
  24'h9e71_c8,
  24'h9e6b_00,
  24'h9e4d_40,
  24'h9e47_2d,
  24'h9e41_6b,
  24'h9e3b_2f,
  24'h9e29_50,
  24'h9e1d_31,
  24'h9e17_35,
  24'h9dcd_0a,
  24'h9dcb_0a,
  24'h9dc9_0a,
  24'h9dae_09,
  24'h9dad_09,
  24'h9dac_09,
  24'h9dab_00,
  24'h9daa_00,
  24'h9da9_00,
  24'h9da8_1e,
  24'h9da7_1e,
  24'h9da6_1e,
  24'h9da5_00,
  24'h9da4_00,
  24'h9da3_00,
  24'h9da2_0f,
  24'h9da1_0f,
  24'h9da0_0f,
  24'h9d9f_1f,
  24'h9d9e_1f,
  24'h9d9d_1f,
  24'h9d9c_3f,
  24'h9d9b_3f,
  24'h9d9a_3f,
  24'h9d99_00,
  24'h9d98_00,
  24'h9d97_00,
  24'h9d96_3f,
  24'h9d95_3f,
  24'h9d94_3f,
  24'h9d83_5a,
  24'h9d7d_42,
  24'h9d75_04,
  24'h9d73_32,
  24'h9d71_c8,
  24'h9d6b_00,
  24'h9d4d_5a,
  24'h9d47_42,
  24'h9d41_6b,
  24'h9d3b_2f,
  24'h9d29_50,
  24'h9d1d_31,
  24'h9d17_35,
  24'h9ccd_0a,
  24'h9ccb_0a,
  24'h9cc9_0a,
  24'h9cc7_40,
  24'h9cc5_40,
  24'h9cc3_40,
  24'h9cc1_50,
  24'h9cbf_50,
  24'h9cbd_50,
  24'h9cae_09,
  24'h9cad_09,
  24'h9cac_09,
  24'h9cab_00,
  24'h9caa_00,
  24'h9ca9_00,
  24'h9ca8_1e,
  24'h9ca7_1e,
  24'h9ca6_1e,
  24'h9ca5_00,
  24'h9ca4_00,
  24'h9ca3_00,
  24'h9ca2_0f,
  24'h9ca1_0f,
  24'h9ca0_0f,
  24'h9c9c_3f,
  24'h9c9b_3f,
  24'h9c9a_3f,
  24'h9c99_00,
  24'h9c98_00,
  24'h9c97_00,
  24'h9c96_3f,
  24'h9c95_3f,
  24'h9c94_3f,
  24'h9c83_40,
  24'h9c7d_2d,
  24'h9c75_04,
  24'h9c73_32,
  24'h9c71_c8,
  24'h9c6b_00,
  24'h9c4d_40,
  24'h9c47_2d,
  24'h9c41_6b,
  24'h9c3b_2f,
  24'h9c29_50,
  24'h9c1d_31,
  24'h9c17_35,
  24'h9a47_00,
  24'h9a46_00,
  24'h9a41_00,
  24'h9a30_05,
  24'h9a2f_05,
  24'h9a2d_03,
  24'h9a2c_01,
  24'h9a27_05,
  24'h9a26_05,
  24'h9a1d_04,
  24'h9a1c_04,
  24'h9a19_00,
  24'h9a14_04,
  24'h9a13_04,
  24'h9955_0a,
  24'h9954_1b,
  24'h9953_8c,
  24'h9952_0a,
  24'h9951_1b,
  24'h9950_8c,
  24'h994f_1b,
  24'h994e_50,
  24'h994d_8c,
  24'h994c_1b,
  24'h994b_50,
  24'h994a_8c,
  24'h9947_3c,
  24'h9944_3c,
  24'h990b_00,
  24'h9909_00,
  24'h9907_00,
  24'h9905_00,
  24'h7b4c_00,
  24'h7b3b_01,
  24'h4421_04,
  24'h3d8a_01,
  24'ha009_c0,
  24'ha007_c0,
  24'ha006_01,
  24'ha005_0a,
  24'ha003_0a,
  24'ha001_0a,
  24'h9a4d_0d,
  24'h9a4c_0d,
  24'h996d_50,
  24'h996c_64,
  24'h996b_8c,
  24'h991a_00,
  24'h9375_64,
  24'h9373_6a,
  24'h9371_6a,
  24'h9205_01,
  24'h9204_71,
  24'h9203_00,
  24'h9202_71,
  24'h9201_6c,
  24'h9200_50,
  24'h9004_03,
  24'h8d27_00,
  24'h8d1f_00,
  24'h7b7d_00,
  24'h7b7c_00,
  24'h7b79_47,
  24'h7b78_0a,
  24'h7b77_08,
  24'h7b76_0b,
  24'h7b75_0e,
  24'h5d77_7f,
  24'h5d38_5a,
  24'h5d37_5a,
  24'h5d26_a8,
  24'h5d25_57,
  24'h5d24_7d,
  24'h5d23_aa,
  24'h5d22_52,
  24'h5d21_0e,
  24'h5d1f_15,
  24'h5d1e_ab,
  24'h5d1d_3a,
  24'h5d1c_45,
  24'h5d1b_a9,
  24'h5d1a_06,
  24'h5d18_8c,
  24'h5d17_65,
  24'h5d16_1d,
  24'h5d15_a3,
  24'h5d14_58,
  24'h5d13_c3,
  24'h5974_01,
  24'h5973_04,
  24'h5757_ff,
  24'h5756_07,
  24'h5755_00,
  24'h5754_00,
  24'h574f_00,
  24'h574e_00,
  24'h574d_ff,
  24'h574c_07,
  24'h55eb_00,
  24'h55ea_00,
  24'h55e9_ff,
  24'h55e8_07,
  24'h55d7_ff,
  24'h55d6_07,
  24'h55d5_00,
  24'h55d4_00,
  24'h38ab_ff,
  24'h38aa_1f,
  24'h38a9_ff,
  24'h38a8_1f,
  24'h4aea_80,
  24'h4ae9_21,
  24'hf61e_04,
  24'hf61c_04,
  24'h4aea_08,
  24'h4ae9_18,
  24'h0808_02,
  24'he07a_01,
  24'he000_00,
  24'h0137_00,
  24'h0136_18,
  24'h0100_00
};

parameter int TOTAL_INIT_OPS = 308;

endpackage
